//-----------------------------------------------------
// Project Name : a.out
// Function     : Execution
// Description  : This is a detailed explanation use several lines to explain everything. You will forget how smart you where when coding this module
// Coder        : G.Cabo
// References   : https://github.com/jaquerinte/MA_2019.git

//***Headers***
`include "defines.vh"
//***Module***
module execute #(
        parameter integer AddrSize = 1
    )
    (
        input  rst_i ,
        input  clk_i ,
        input  wreg_i ,
        input  m2reg_i ,
        input  wmem_i ,
        input  aluc_i ,
        input  aluimm_i ,
        input  [`BITS_REGFILE : 0] destination_i ,
        input  [AddrSize - 1 : 0] op1_i ,
        input  [AddrSize - 1 : 0] op2_i ,
        input  [AddrSize - 1 : 0] extendedimm_i ,
        output wreg_o ,
        output m2reg_o ,
        output wmem_o ,
        output [`BITS_REGFILE : 0] destination_o ,
        output [AddrSize - 1 : 0] aluresult_o ,
        output [AddrSize - 1 : 0] op2_o 
    );



//***Interal logic generated by compiler***  
//***Handcrafted Internal logic*** 
//TODO
endmodule
