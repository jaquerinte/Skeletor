//-----------------------------------------------------
// Project Name : a.out

//***Headers***
//***Module***
module decode #(
        parameter integer AddrSize = 1,
        parameter integer BITS_REGFILE = 1
    )
    (
        input  clk_i ,
        input  rst_i ,
        input  [AddrSize - 1 : 0] instruction_i ,
        input  [BITS_REGFILE - 1 : 0] destination_i ,
        input  [AddrSize - 1 : 0] datareg_i ,
        input  wreg_i ,
        output wreg_o ,
        output m2reg_o ,
        output wmem_o ,
        output aluc_o ,
        output aluimm_o ,
        output [BITS_REGFILE : 0] destination_o ,
        output [AddrSize - 1 : 0] op1_o ,
        output [AddrSize - 1 : 0] op2_o ,
        output [AddrSize - 1 : 0] extendedimm_o 
    );

//***Interal logic generated by compiler***  


//***Handcrafted Internal logic*** 
//TODO
endmodule
