//-------------------------------------------------
// Generated defines from vericon
//-------------------------------------------------

`define ADDR_SIZE 32 
`define T_ADDR_SIZE 32 

