//-----------------------------------------------------
// Project Name : a.out
// Function     : Decode instructions and operand fetch
// Description  : This is a detailed explanation use several lines to explain everything. You will forget how smart you where when coding this module
// Coder        : G.Cabo
// References   : https://github.com/jaquerinte/MA_2019.git

//***Headers***
`include "defines.vh"
//***Module***
module decode #(
        parameter integer AddrSize = 1
    )
    (
        input  rst_i ,
        input  clk_i ,
        input  [AddrSize - 1 : 0] instruction_i ,
        input  [`BITS_REGFILE - 1 : 0] destination_i ,
        input  [AddrSize - 1 : 0] datareg_i ,
        input  wreg_i ,
        output wreg_o ,
        output m2reg_o ,
        output wmem_o ,
        output aluc_o ,
        output aluimm_o ,
        output [`BITS_REGFILE : 0] destination_o ,
        output [AddrSize - 1 : 0] op1_o ,
        output [AddrSize - 1 : 0] op2_o ,
        output [AddrSize - 1 : 0] extendedimm_o 
    );



//***Interal logic generated by compiler***  
//***Handcrafted Internal logic*** 
//TODO
endmodule
