//-----------------------------------------------------
// Project Name : a.out
// Function     : Fetch instructions
// Description  : This is a detailed explanation use several lines to explain everything. You will forget how smart you where when coding this module
// Coder        : G.Cabo
// References   : https://github.com/jaquerinte/MA_2019.git

//***Headers***
`include "defines.vh"
//***Module***
module fetch #(
        parameter integer AddrSize = 1
    )
    (
        input  rst_i ,
        input  clk_i ,
        input  [AddrSize - 1 : 0] pc_i ,
        output [AddrSize - 1 : 0] nextpc_o ,
        output [AddrSize - 1 : 0] instruction_o 
    );



//***Interal logic generated by compiler***  
//***Handcrafted Internal logic*** 
//TODO
endmodule
