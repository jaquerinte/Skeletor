//-----------------------------------------------------
// Project Name : a.out

//***Headers***
//***Module***
module writeback #(
        parameter integer AddrSize = 1,
        parameter integer BITS_REGFILE = 1
    )
    (
        input  clk_i ,
        input  rst_i ,
        input  wreg_i ,
        input  m2reg_i ,
        input  [AddrSize - 1 : 0] aluresult_i ,
        input  [AddrSize - 1 : 0] dmemout_i ,
        input  [BITS_REGFILE : 0] destination_i ,
        output wreg_o ,
        output [BITS_REGFILE : 0] destination_o ,
        output [AddrSize - 1 : 0] datareg_o 
    );

//***Interal logic generated by compiler***  


//***Handcrafted Internal logic*** 
//TODO
endmodule
