//-------------------------------------------------
// Generated defines                               
//-------------------------------------------------

`define ADDR_SIZE 32
`define BITS_REGFILE 5
//-------------------------------------------------
// Generated defines                               
//-------------------------------------------------

`define ADDR_SIZE 32
`define BITS_REGFILE 5
//-------------------------------------------------
// Generated defines                               
//-------------------------------------------------

`define ADDR_SIZE 32
`define BITS_REGFILE 5
//-------------------------------------------------
// Generated defines                               
//-------------------------------------------------

`define ADDR_SIZE 32
`define BITS_REGFILE 5
//-------------------------------------------------
// Generated defines                               
//-------------------------------------------------

`define ADDR_SIZE 32
`define BITS_REGFILE 5
//-------------------------------------------------
// Generated defines                               
//-------------------------------------------------

`define ADDR_SIZE 32
`define BITS_REGFILE 5
