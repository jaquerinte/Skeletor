//-----------------------------------------------------
// Project Name : Sample_Code
// File Name    : Module name
// Function     : rdy_o is high when a n bit counter overflow 
// Description  : This is a detailed explanation use several
//                lines to explain everything. You will forget
//                how smart you where when coding this module
// Coder        : G.Cabo
// References   : https://github.com/jaquerinte/MA_2019.git
//-----------------------------------------------------

//***Headers***
//***Module***
module c #(
        parameter integer n  = 2    //Size of counter 
    )
    (
        input rst_i,    //Reset when high connected to top
        input clk_i,    //Clock generated by top
        output rdy_o    //Ready generated by A
    );
    //***Interal logic generated by compiler***  
    //***Handcrafted Internal logic*** 
    //TODO: This module has a n bits counter that triggers rdy_o at overflow
    reg rdy_int;
    assign rdy_o = rdy_int; 
    
    reg [n-1:0] value;
    always@(posedge clk_i) begin
        if(rst_i)
            value<=0;
        else begin
            value<=value+1;
            if({n{1'b0}} == ~value)//if all bits are 1 then overflow
                rdy_int<=1;
            else
                rdy_int<=0;
        end
    end 
endmodule

